LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Generic_MUX_4to1 is
	GENERIC
	(
		N	:	INTEGER
	);
	
	PORT
	(
		IN_A	:	IN		STD_LOGIC_VECTOR	(N-1 DOWNTO 0);
		IN_B	:	IN		STD_LOGIC_VECTOR	(N-1 DOWNTO 0);
		IN_C	:	IN		STD_LOGIC_VECTOR	(N-1 DOWNTO 0);
		IN_D	:	IN		STD_LOGIC_VECTOR	(N-1 DOWNTO 0);
		OUT_X	:	OUT	STD_LOGIC_VECTOR	(N-1 DOWNTO 0);
		SEL	:	IN		STD_LOGIC_VECTOR	(1   DOWNTO 0)
	);
END Generic_MUX_4to1;

ARCHITECTURE Gen_MUX_4to1 OF Generic_MUX_4to1 IS
BEGIN
	Generic_MUX_4_to_1 : PROCESS(IN_A,IN_B,IN_C,IN_D,SEL)
	BEGIN
		CASE SEL IS
			WHEN "00"	=>	OUT_X	<= IN_A;
			WHEN "01"	=>	OUT_X	<= IN_B;
			WHEN "10"	=>	OUT_X	<= IN_C;
			WHEN OTHERS	=>	OUT_X	<= IN_D;
		END CASE;
	END PROCESS Generic_MUX_4_to_1;
END Gen_MUX_4to1;