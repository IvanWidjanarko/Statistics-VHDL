LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Generic_MUX_2to1 is
	GENERIC
	(
		N	:	INTEGER
	);
	
	PORT
	(
		IN_A	:	IN		STD_LOGIC_VECTOR	(N-1 DOWNTO 0);
		IN_B	:	IN		STD_LOGIC_VECTOR	(N-1 DOWNTO 0);
		OUT_X	:	OUT	STD_LOGIC_VECTOR	(N-1 DOWNTO 0);
		SEL	:	IN		STD_LOGIC
	);
END Generic_MUX_2to1;

ARCHITECTURE Gen_MUX_2to1 OF Generic_MUX_2to1 IS
BEGIN
	Generic_MUX_2_to_1 : PROCESS(IN_A,IN_B,SEL)
	BEGIN
		IF SEL = '0' THEN
			OUT_X <= IN_A;
		ELSE
			OUT_X <= IN_B;
		END IF;
	END PROCESS Generic_MUX_2_to_1;
END Gen_MUX_2to1;